`timescale 1ns/1ps

module radix2_tb ();
	/****************************************************************************
    * Parameter
    ***************************************************************************/
	parameter WIDTH = 18;
	parameter psi = 3383;

   /****************************************************************************
    * Signals
    ***************************************************************************/

   reg signed [WIDTH-1:0] in1;
   reg signed [WIDTH-1:0] in2;
   reg signed [WIDTH-1:0] w1;
   reg signed [WIDTH-1:0] w2;
   wire signed[WIDTH-1:0] out1;
   wire signed[WIDTH-1:0] out2;

   /****************************************************************************
    * Generate Clock Signals
    ***************************************************************************/

   /****************************************************************************
    * Instantiate Modules
    ***************************************************************************/

   Radix_2 #(.WIDTH(WIDTH)) uut (
      .input_1		(in1),
		.input_2		(in2),
		.weight_1	(w1),
		.weight_2	(w2),
		.output_1	(out1),
		.output_2	(out2)
   );

   /****************************************************************************
    * Apply Stimulus
    ***************************************************************************/

   initial begin
		$dumpfile("wave.vcd");
		$dumpvars(0,radix2_tb);

		in1 = 1;
		in2 = 2;
		w1 = 1;
		w2 = 256;
		#1;
		$display ("Result 1: %b (%d) ", out1, out1);
		$display ("Result 2: %b (%d) ", out2, out2);

		
      $finish;

   end

endmodule
