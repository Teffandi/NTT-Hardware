parameter width = 32,
parameter w1= 1,
parameter w2= 1925,
parameter w3= 3383,
parameter w4= 6468