`timescale 1ns/1ps

module modulo_tb ();
	/****************************************************************************
    * Parameter
    ***************************************************************************/
	parameter width = 18;
	parameter m = 16;

   /****************************************************************************
    * Signals
    ***************************************************************************/

   reg signed [2*m+2:0] in;
   wire [width-1:0] out;

   /****************************************************************************
    * Generate Clock Signals
    ***************************************************************************/


   /****************************************************************************
    * Instantiate Modules
    ***************************************************************************/

   modulo #(.WIDTH(width), .m(m)) uut (
      .input_mod		(in),
      .output_mod  	(out)
   );

   /****************************************************************************
    * Apply Stimulus
    ***************************************************************************/

   initial begin
		$dumpfile("wave.vcd");
		$dumpvars(0,modulo_tb);

		in = 0;
		#1;
		$display ("%b (%d) mod 65537 = %b (%d)", in, in, out, out);

		in = 65537;
		#1;
		$display ("%b (%d) mod 65537 = %b (%d)", in, in, out, out);

		in = 65540;
		#1;
		$display ("%b (%d) mod 65537 = %b (%d)", in, in, out, out);

		in = -1;
		#1;
		$display ("%b (%d) mod 65537 = %b (%d)", in, in, out, out);

		in = -48577;
		#1;
		$display ("%b (%d) mod 65537 = %b (%d)", in, in, out, out);

      $finish;

   end

endmodule
