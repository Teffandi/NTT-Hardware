parameter width = 32