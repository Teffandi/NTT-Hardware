parameter width = 16